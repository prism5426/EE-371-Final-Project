module game_logic(clk, resetGame, press, x, y, r, g, b);
	 input logic clk, resetGame, press;
    input logic [9:0] x;
    input logic [8:0] y;
    output logic [7:0] r, g, b;
	

endmodule
